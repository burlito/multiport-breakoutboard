.title KiCad schematic
SW1 /GND Net-_R1-Pad1_ /33V SW_SPDT_MSM
J4 /PWR_TGL /GND /VID_OUT /AUDIO_L /AUDIO_R /SLCT /RX /TX /XRST /33V MULT_terminal
R1 Net-_R1-Pad1_ /SLCT 100R
J1 /VBUS /USB_D- /USB_D+ /USB_ID /USB_GND USB_terminal
J2 /VBUS /USB_D- /USB_D+ /USB_ID /USB_GND /USB_GND USB_B_Micro
J3 /PWR_TGL /GND /VID_OUT /AUDIO_L /AUDIO_R /SLCT /RX /TX /XRST /33V /USB_GND /USB_ID /USB_D+ /USB_D- /VBUS soldier_pads
.end
